// FETCH
//

module fetcher (
input logic clk, reset, enable, zero,
output logic c_out, zero_out
);



endmodule