//RAM
module RAM();

endmodule 