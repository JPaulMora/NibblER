module busDriver(
    input enable;
    
)