module In(
    input [3:0] A,
    inout [3:0] Y
);

assign Y = ()
