//PC COUNTER

module pcCounter(clk, reset, incPC, loadPC, outValue, loadValues);
    output [11:0] outValue, loadValues;
    input clk, reset, loadPC, incPC;
    
endmodule